library verilog;
use verilog.vl_types.all;
entity vending_machine_vlg_vec_tst is
end vending_machine_vlg_vec_tst;
