library verilog;
use verilog.vl_types.all;
entity acumulador8_vlg_vec_tst is
end acumulador8_vlg_vec_tst;
